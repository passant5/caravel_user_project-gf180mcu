magic
tech gf180mcuC
magscale 1 5
timestamp 1670786345
<< obsm1 >>
rect 672 1079 89320 58438
<< metal2 >>
rect 672 59600 728 60000
rect 1456 59600 1512 60000
rect 2240 59600 2296 60000
rect 3024 59600 3080 60000
rect 3808 59600 3864 60000
rect 4592 59600 4648 60000
rect 5376 59600 5432 60000
rect 6160 59600 6216 60000
rect 6944 59600 7000 60000
rect 7728 59600 7784 60000
rect 8512 59600 8568 60000
rect 9296 59600 9352 60000
rect 10080 59600 10136 60000
rect 10864 59600 10920 60000
rect 11648 59600 11704 60000
rect 12432 59600 12488 60000
rect 13216 59600 13272 60000
rect 14000 59600 14056 60000
rect 14784 59600 14840 60000
rect 15568 59600 15624 60000
rect 16352 59600 16408 60000
rect 17136 59600 17192 60000
rect 17920 59600 17976 60000
rect 18704 59600 18760 60000
rect 19488 59600 19544 60000
rect 20272 59600 20328 60000
rect 21056 59600 21112 60000
rect 21840 59600 21896 60000
rect 22624 59600 22680 60000
rect 23408 59600 23464 60000
rect 24192 59600 24248 60000
rect 24976 59600 25032 60000
rect 25760 59600 25816 60000
rect 26544 59600 26600 60000
rect 27328 59600 27384 60000
rect 28112 59600 28168 60000
rect 28896 59600 28952 60000
rect 29680 59600 29736 60000
rect 30464 59600 30520 60000
rect 31248 59600 31304 60000
rect 32032 59600 32088 60000
rect 32816 59600 32872 60000
rect 33600 59600 33656 60000
rect 34384 59600 34440 60000
rect 35168 59600 35224 60000
rect 35952 59600 36008 60000
rect 36736 59600 36792 60000
rect 37520 59600 37576 60000
rect 38304 59600 38360 60000
rect 39088 59600 39144 60000
rect 39872 59600 39928 60000
rect 40656 59600 40712 60000
rect 41440 59600 41496 60000
rect 42224 59600 42280 60000
rect 43008 59600 43064 60000
rect 43792 59600 43848 60000
rect 44576 59600 44632 60000
rect 45360 59600 45416 60000
rect 46144 59600 46200 60000
rect 46928 59600 46984 60000
rect 47712 59600 47768 60000
rect 48496 59600 48552 60000
rect 49280 59600 49336 60000
rect 50064 59600 50120 60000
rect 50848 59600 50904 60000
rect 51632 59600 51688 60000
rect 52416 59600 52472 60000
rect 53200 59600 53256 60000
rect 53984 59600 54040 60000
rect 54768 59600 54824 60000
rect 55552 59600 55608 60000
rect 56336 59600 56392 60000
rect 57120 59600 57176 60000
rect 57904 59600 57960 60000
rect 58688 59600 58744 60000
rect 59472 59600 59528 60000
rect 60256 59600 60312 60000
rect 61040 59600 61096 60000
rect 61824 59600 61880 60000
rect 62608 59600 62664 60000
rect 63392 59600 63448 60000
rect 64176 59600 64232 60000
rect 64960 59600 65016 60000
rect 65744 59600 65800 60000
rect 66528 59600 66584 60000
rect 67312 59600 67368 60000
rect 68096 59600 68152 60000
rect 68880 59600 68936 60000
rect 69664 59600 69720 60000
rect 70448 59600 70504 60000
rect 71232 59600 71288 60000
rect 72016 59600 72072 60000
rect 72800 59600 72856 60000
rect 73584 59600 73640 60000
rect 74368 59600 74424 60000
rect 75152 59600 75208 60000
rect 75936 59600 75992 60000
rect 76720 59600 76776 60000
rect 77504 59600 77560 60000
rect 78288 59600 78344 60000
rect 79072 59600 79128 60000
rect 79856 59600 79912 60000
rect 80640 59600 80696 60000
rect 81424 59600 81480 60000
rect 82208 59600 82264 60000
rect 82992 59600 83048 60000
rect 83776 59600 83832 60000
rect 84560 59600 84616 60000
rect 85344 59600 85400 60000
rect 86128 59600 86184 60000
rect 86912 59600 86968 60000
rect 87696 59600 87752 60000
rect 88480 59600 88536 60000
rect 89264 59600 89320 60000
rect 2800 0 2856 400
rect 3080 0 3136 400
rect 3360 0 3416 400
rect 3640 0 3696 400
rect 3920 0 3976 400
rect 4200 0 4256 400
rect 4480 0 4536 400
rect 4760 0 4816 400
rect 5040 0 5096 400
rect 5320 0 5376 400
rect 5600 0 5656 400
rect 5880 0 5936 400
rect 6160 0 6216 400
rect 6440 0 6496 400
rect 6720 0 6776 400
rect 7000 0 7056 400
rect 7280 0 7336 400
rect 7560 0 7616 400
rect 7840 0 7896 400
rect 8120 0 8176 400
rect 8400 0 8456 400
rect 8680 0 8736 400
rect 8960 0 9016 400
rect 9240 0 9296 400
rect 9520 0 9576 400
rect 9800 0 9856 400
rect 10080 0 10136 400
rect 10360 0 10416 400
rect 10640 0 10696 400
rect 10920 0 10976 400
rect 11200 0 11256 400
rect 11480 0 11536 400
rect 11760 0 11816 400
rect 12040 0 12096 400
rect 12320 0 12376 400
rect 12600 0 12656 400
rect 12880 0 12936 400
rect 13160 0 13216 400
rect 13440 0 13496 400
rect 13720 0 13776 400
rect 14000 0 14056 400
rect 14280 0 14336 400
rect 14560 0 14616 400
rect 14840 0 14896 400
rect 15120 0 15176 400
rect 15400 0 15456 400
rect 15680 0 15736 400
rect 15960 0 16016 400
rect 16240 0 16296 400
rect 16520 0 16576 400
rect 16800 0 16856 400
rect 17080 0 17136 400
rect 17360 0 17416 400
rect 17640 0 17696 400
rect 17920 0 17976 400
rect 18200 0 18256 400
rect 18480 0 18536 400
rect 18760 0 18816 400
rect 19040 0 19096 400
rect 19320 0 19376 400
rect 19600 0 19656 400
rect 19880 0 19936 400
rect 20160 0 20216 400
rect 20440 0 20496 400
rect 20720 0 20776 400
rect 21000 0 21056 400
rect 21280 0 21336 400
rect 21560 0 21616 400
rect 21840 0 21896 400
rect 22120 0 22176 400
rect 22400 0 22456 400
rect 22680 0 22736 400
rect 22960 0 23016 400
rect 23240 0 23296 400
rect 23520 0 23576 400
rect 23800 0 23856 400
rect 24080 0 24136 400
rect 24360 0 24416 400
rect 24640 0 24696 400
rect 24920 0 24976 400
rect 25200 0 25256 400
rect 25480 0 25536 400
rect 25760 0 25816 400
rect 26040 0 26096 400
rect 26320 0 26376 400
rect 26600 0 26656 400
rect 26880 0 26936 400
rect 27160 0 27216 400
rect 27440 0 27496 400
rect 27720 0 27776 400
rect 28000 0 28056 400
rect 28280 0 28336 400
rect 28560 0 28616 400
rect 28840 0 28896 400
rect 29120 0 29176 400
rect 29400 0 29456 400
rect 29680 0 29736 400
rect 29960 0 30016 400
rect 30240 0 30296 400
rect 30520 0 30576 400
rect 30800 0 30856 400
rect 31080 0 31136 400
rect 31360 0 31416 400
rect 31640 0 31696 400
rect 31920 0 31976 400
rect 32200 0 32256 400
rect 32480 0 32536 400
rect 32760 0 32816 400
rect 33040 0 33096 400
rect 33320 0 33376 400
rect 33600 0 33656 400
rect 33880 0 33936 400
rect 34160 0 34216 400
rect 34440 0 34496 400
rect 34720 0 34776 400
rect 35000 0 35056 400
rect 35280 0 35336 400
rect 35560 0 35616 400
rect 35840 0 35896 400
rect 36120 0 36176 400
rect 36400 0 36456 400
rect 36680 0 36736 400
rect 36960 0 37016 400
rect 37240 0 37296 400
rect 37520 0 37576 400
rect 37800 0 37856 400
rect 38080 0 38136 400
rect 38360 0 38416 400
rect 38640 0 38696 400
rect 38920 0 38976 400
rect 39200 0 39256 400
rect 39480 0 39536 400
rect 39760 0 39816 400
rect 40040 0 40096 400
rect 40320 0 40376 400
rect 40600 0 40656 400
rect 40880 0 40936 400
rect 41160 0 41216 400
rect 41440 0 41496 400
rect 41720 0 41776 400
rect 42000 0 42056 400
rect 42280 0 42336 400
rect 42560 0 42616 400
rect 42840 0 42896 400
rect 43120 0 43176 400
rect 43400 0 43456 400
rect 43680 0 43736 400
rect 43960 0 44016 400
rect 44240 0 44296 400
rect 44520 0 44576 400
rect 44800 0 44856 400
rect 45080 0 45136 400
rect 45360 0 45416 400
rect 45640 0 45696 400
rect 45920 0 45976 400
rect 46200 0 46256 400
rect 46480 0 46536 400
rect 46760 0 46816 400
rect 47040 0 47096 400
rect 47320 0 47376 400
rect 47600 0 47656 400
rect 47880 0 47936 400
rect 48160 0 48216 400
rect 48440 0 48496 400
rect 48720 0 48776 400
rect 49000 0 49056 400
rect 49280 0 49336 400
rect 49560 0 49616 400
rect 49840 0 49896 400
rect 50120 0 50176 400
rect 50400 0 50456 400
rect 50680 0 50736 400
rect 50960 0 51016 400
rect 51240 0 51296 400
rect 51520 0 51576 400
rect 51800 0 51856 400
rect 52080 0 52136 400
rect 52360 0 52416 400
rect 52640 0 52696 400
rect 52920 0 52976 400
rect 53200 0 53256 400
rect 53480 0 53536 400
rect 53760 0 53816 400
rect 54040 0 54096 400
rect 54320 0 54376 400
rect 54600 0 54656 400
rect 54880 0 54936 400
rect 55160 0 55216 400
rect 55440 0 55496 400
rect 55720 0 55776 400
rect 56000 0 56056 400
rect 56280 0 56336 400
rect 56560 0 56616 400
rect 56840 0 56896 400
rect 57120 0 57176 400
rect 57400 0 57456 400
rect 57680 0 57736 400
rect 57960 0 58016 400
rect 58240 0 58296 400
rect 58520 0 58576 400
rect 58800 0 58856 400
rect 59080 0 59136 400
rect 59360 0 59416 400
rect 59640 0 59696 400
rect 59920 0 59976 400
rect 60200 0 60256 400
rect 60480 0 60536 400
rect 60760 0 60816 400
rect 61040 0 61096 400
rect 61320 0 61376 400
rect 61600 0 61656 400
rect 61880 0 61936 400
rect 62160 0 62216 400
rect 62440 0 62496 400
rect 62720 0 62776 400
rect 63000 0 63056 400
rect 63280 0 63336 400
rect 63560 0 63616 400
rect 63840 0 63896 400
rect 64120 0 64176 400
rect 64400 0 64456 400
rect 64680 0 64736 400
rect 64960 0 65016 400
rect 65240 0 65296 400
rect 65520 0 65576 400
rect 65800 0 65856 400
rect 66080 0 66136 400
rect 66360 0 66416 400
rect 66640 0 66696 400
rect 66920 0 66976 400
rect 67200 0 67256 400
rect 67480 0 67536 400
rect 67760 0 67816 400
rect 68040 0 68096 400
rect 68320 0 68376 400
rect 68600 0 68656 400
rect 68880 0 68936 400
rect 69160 0 69216 400
rect 69440 0 69496 400
rect 69720 0 69776 400
rect 70000 0 70056 400
rect 70280 0 70336 400
rect 70560 0 70616 400
rect 70840 0 70896 400
rect 71120 0 71176 400
rect 71400 0 71456 400
rect 71680 0 71736 400
rect 71960 0 72016 400
rect 72240 0 72296 400
rect 72520 0 72576 400
rect 72800 0 72856 400
rect 73080 0 73136 400
rect 73360 0 73416 400
rect 73640 0 73696 400
rect 73920 0 73976 400
rect 74200 0 74256 400
rect 74480 0 74536 400
rect 74760 0 74816 400
rect 75040 0 75096 400
rect 75320 0 75376 400
rect 75600 0 75656 400
rect 75880 0 75936 400
rect 76160 0 76216 400
rect 76440 0 76496 400
rect 76720 0 76776 400
rect 77000 0 77056 400
rect 77280 0 77336 400
rect 77560 0 77616 400
rect 77840 0 77896 400
rect 78120 0 78176 400
rect 78400 0 78456 400
rect 78680 0 78736 400
rect 78960 0 79016 400
rect 79240 0 79296 400
rect 79520 0 79576 400
rect 79800 0 79856 400
rect 80080 0 80136 400
rect 80360 0 80416 400
rect 80640 0 80696 400
rect 80920 0 80976 400
rect 81200 0 81256 400
rect 81480 0 81536 400
rect 81760 0 81816 400
rect 82040 0 82096 400
rect 82320 0 82376 400
rect 82600 0 82656 400
rect 82880 0 82936 400
rect 83160 0 83216 400
rect 83440 0 83496 400
rect 83720 0 83776 400
rect 84000 0 84056 400
rect 84280 0 84336 400
rect 84560 0 84616 400
rect 84840 0 84896 400
rect 85120 0 85176 400
rect 85400 0 85456 400
rect 85680 0 85736 400
rect 85960 0 86016 400
rect 86240 0 86296 400
rect 86520 0 86576 400
rect 86800 0 86856 400
rect 87080 0 87136 400
<< obsm2 >>
rect 14 59570 642 59682
rect 758 59570 1426 59682
rect 1542 59570 2210 59682
rect 2326 59570 2994 59682
rect 3110 59570 3778 59682
rect 3894 59570 4562 59682
rect 4678 59570 5346 59682
rect 5462 59570 6130 59682
rect 6246 59570 6914 59682
rect 7030 59570 7698 59682
rect 7814 59570 8482 59682
rect 8598 59570 9266 59682
rect 9382 59570 10050 59682
rect 10166 59570 10834 59682
rect 10950 59570 11618 59682
rect 11734 59570 12402 59682
rect 12518 59570 13186 59682
rect 13302 59570 13970 59682
rect 14086 59570 14754 59682
rect 14870 59570 15538 59682
rect 15654 59570 16322 59682
rect 16438 59570 17106 59682
rect 17222 59570 17890 59682
rect 18006 59570 18674 59682
rect 18790 59570 19458 59682
rect 19574 59570 20242 59682
rect 20358 59570 21026 59682
rect 21142 59570 21810 59682
rect 21926 59570 22594 59682
rect 22710 59570 23378 59682
rect 23494 59570 24162 59682
rect 24278 59570 24946 59682
rect 25062 59570 25730 59682
rect 25846 59570 26514 59682
rect 26630 59570 27298 59682
rect 27414 59570 28082 59682
rect 28198 59570 28866 59682
rect 28982 59570 29650 59682
rect 29766 59570 30434 59682
rect 30550 59570 31218 59682
rect 31334 59570 32002 59682
rect 32118 59570 32786 59682
rect 32902 59570 33570 59682
rect 33686 59570 34354 59682
rect 34470 59570 35138 59682
rect 35254 59570 35922 59682
rect 36038 59570 36706 59682
rect 36822 59570 37490 59682
rect 37606 59570 38274 59682
rect 38390 59570 39058 59682
rect 39174 59570 39842 59682
rect 39958 59570 40626 59682
rect 40742 59570 41410 59682
rect 41526 59570 42194 59682
rect 42310 59570 42978 59682
rect 43094 59570 43762 59682
rect 43878 59570 44546 59682
rect 44662 59570 45330 59682
rect 45446 59570 46114 59682
rect 46230 59570 46898 59682
rect 47014 59570 47682 59682
rect 47798 59570 48466 59682
rect 48582 59570 49250 59682
rect 49366 59570 50034 59682
rect 50150 59570 50818 59682
rect 50934 59570 51602 59682
rect 51718 59570 52386 59682
rect 52502 59570 53170 59682
rect 53286 59570 53954 59682
rect 54070 59570 54738 59682
rect 54854 59570 55522 59682
rect 55638 59570 56306 59682
rect 56422 59570 57090 59682
rect 57206 59570 57874 59682
rect 57990 59570 58658 59682
rect 58774 59570 59442 59682
rect 59558 59570 60226 59682
rect 60342 59570 61010 59682
rect 61126 59570 61794 59682
rect 61910 59570 62578 59682
rect 62694 59570 63362 59682
rect 63478 59570 64146 59682
rect 64262 59570 64930 59682
rect 65046 59570 65714 59682
rect 65830 59570 66498 59682
rect 66614 59570 67282 59682
rect 67398 59570 68066 59682
rect 68182 59570 68850 59682
rect 68966 59570 69634 59682
rect 69750 59570 70418 59682
rect 70534 59570 71202 59682
rect 71318 59570 71986 59682
rect 72102 59570 72770 59682
rect 72886 59570 73554 59682
rect 73670 59570 74338 59682
rect 74454 59570 75122 59682
rect 75238 59570 75906 59682
rect 76022 59570 76690 59682
rect 76806 59570 77474 59682
rect 77590 59570 78258 59682
rect 78374 59570 79042 59682
rect 79158 59570 79826 59682
rect 79942 59570 80610 59682
rect 80726 59570 81394 59682
rect 81510 59570 82178 59682
rect 82294 59570 82962 59682
rect 83078 59570 83746 59682
rect 83862 59570 84530 59682
rect 84646 59570 85314 59682
rect 85430 59570 86098 59682
rect 86214 59570 86882 59682
rect 86998 59570 87666 59682
rect 87782 59570 88450 59682
rect 88566 59570 89234 59682
rect 14 430 89306 59570
rect 14 400 2770 430
rect 2886 400 3050 430
rect 3166 400 3330 430
rect 3446 400 3610 430
rect 3726 400 3890 430
rect 4006 400 4170 430
rect 4286 400 4450 430
rect 4566 400 4730 430
rect 4846 400 5010 430
rect 5126 400 5290 430
rect 5406 400 5570 430
rect 5686 400 5850 430
rect 5966 400 6130 430
rect 6246 400 6410 430
rect 6526 400 6690 430
rect 6806 400 6970 430
rect 7086 400 7250 430
rect 7366 400 7530 430
rect 7646 400 7810 430
rect 7926 400 8090 430
rect 8206 400 8370 430
rect 8486 400 8650 430
rect 8766 400 8930 430
rect 9046 400 9210 430
rect 9326 400 9490 430
rect 9606 400 9770 430
rect 9886 400 10050 430
rect 10166 400 10330 430
rect 10446 400 10610 430
rect 10726 400 10890 430
rect 11006 400 11170 430
rect 11286 400 11450 430
rect 11566 400 11730 430
rect 11846 400 12010 430
rect 12126 400 12290 430
rect 12406 400 12570 430
rect 12686 400 12850 430
rect 12966 400 13130 430
rect 13246 400 13410 430
rect 13526 400 13690 430
rect 13806 400 13970 430
rect 14086 400 14250 430
rect 14366 400 14530 430
rect 14646 400 14810 430
rect 14926 400 15090 430
rect 15206 400 15370 430
rect 15486 400 15650 430
rect 15766 400 15930 430
rect 16046 400 16210 430
rect 16326 400 16490 430
rect 16606 400 16770 430
rect 16886 400 17050 430
rect 17166 400 17330 430
rect 17446 400 17610 430
rect 17726 400 17890 430
rect 18006 400 18170 430
rect 18286 400 18450 430
rect 18566 400 18730 430
rect 18846 400 19010 430
rect 19126 400 19290 430
rect 19406 400 19570 430
rect 19686 400 19850 430
rect 19966 400 20130 430
rect 20246 400 20410 430
rect 20526 400 20690 430
rect 20806 400 20970 430
rect 21086 400 21250 430
rect 21366 400 21530 430
rect 21646 400 21810 430
rect 21926 400 22090 430
rect 22206 400 22370 430
rect 22486 400 22650 430
rect 22766 400 22930 430
rect 23046 400 23210 430
rect 23326 400 23490 430
rect 23606 400 23770 430
rect 23886 400 24050 430
rect 24166 400 24330 430
rect 24446 400 24610 430
rect 24726 400 24890 430
rect 25006 400 25170 430
rect 25286 400 25450 430
rect 25566 400 25730 430
rect 25846 400 26010 430
rect 26126 400 26290 430
rect 26406 400 26570 430
rect 26686 400 26850 430
rect 26966 400 27130 430
rect 27246 400 27410 430
rect 27526 400 27690 430
rect 27806 400 27970 430
rect 28086 400 28250 430
rect 28366 400 28530 430
rect 28646 400 28810 430
rect 28926 400 29090 430
rect 29206 400 29370 430
rect 29486 400 29650 430
rect 29766 400 29930 430
rect 30046 400 30210 430
rect 30326 400 30490 430
rect 30606 400 30770 430
rect 30886 400 31050 430
rect 31166 400 31330 430
rect 31446 400 31610 430
rect 31726 400 31890 430
rect 32006 400 32170 430
rect 32286 400 32450 430
rect 32566 400 32730 430
rect 32846 400 33010 430
rect 33126 400 33290 430
rect 33406 400 33570 430
rect 33686 400 33850 430
rect 33966 400 34130 430
rect 34246 400 34410 430
rect 34526 400 34690 430
rect 34806 400 34970 430
rect 35086 400 35250 430
rect 35366 400 35530 430
rect 35646 400 35810 430
rect 35926 400 36090 430
rect 36206 400 36370 430
rect 36486 400 36650 430
rect 36766 400 36930 430
rect 37046 400 37210 430
rect 37326 400 37490 430
rect 37606 400 37770 430
rect 37886 400 38050 430
rect 38166 400 38330 430
rect 38446 400 38610 430
rect 38726 400 38890 430
rect 39006 400 39170 430
rect 39286 400 39450 430
rect 39566 400 39730 430
rect 39846 400 40010 430
rect 40126 400 40290 430
rect 40406 400 40570 430
rect 40686 400 40850 430
rect 40966 400 41130 430
rect 41246 400 41410 430
rect 41526 400 41690 430
rect 41806 400 41970 430
rect 42086 400 42250 430
rect 42366 400 42530 430
rect 42646 400 42810 430
rect 42926 400 43090 430
rect 43206 400 43370 430
rect 43486 400 43650 430
rect 43766 400 43930 430
rect 44046 400 44210 430
rect 44326 400 44490 430
rect 44606 400 44770 430
rect 44886 400 45050 430
rect 45166 400 45330 430
rect 45446 400 45610 430
rect 45726 400 45890 430
rect 46006 400 46170 430
rect 46286 400 46450 430
rect 46566 400 46730 430
rect 46846 400 47010 430
rect 47126 400 47290 430
rect 47406 400 47570 430
rect 47686 400 47850 430
rect 47966 400 48130 430
rect 48246 400 48410 430
rect 48526 400 48690 430
rect 48806 400 48970 430
rect 49086 400 49250 430
rect 49366 400 49530 430
rect 49646 400 49810 430
rect 49926 400 50090 430
rect 50206 400 50370 430
rect 50486 400 50650 430
rect 50766 400 50930 430
rect 51046 400 51210 430
rect 51326 400 51490 430
rect 51606 400 51770 430
rect 51886 400 52050 430
rect 52166 400 52330 430
rect 52446 400 52610 430
rect 52726 400 52890 430
rect 53006 400 53170 430
rect 53286 400 53450 430
rect 53566 400 53730 430
rect 53846 400 54010 430
rect 54126 400 54290 430
rect 54406 400 54570 430
rect 54686 400 54850 430
rect 54966 400 55130 430
rect 55246 400 55410 430
rect 55526 400 55690 430
rect 55806 400 55970 430
rect 56086 400 56250 430
rect 56366 400 56530 430
rect 56646 400 56810 430
rect 56926 400 57090 430
rect 57206 400 57370 430
rect 57486 400 57650 430
rect 57766 400 57930 430
rect 58046 400 58210 430
rect 58326 400 58490 430
rect 58606 400 58770 430
rect 58886 400 59050 430
rect 59166 400 59330 430
rect 59446 400 59610 430
rect 59726 400 59890 430
rect 60006 400 60170 430
rect 60286 400 60450 430
rect 60566 400 60730 430
rect 60846 400 61010 430
rect 61126 400 61290 430
rect 61406 400 61570 430
rect 61686 400 61850 430
rect 61966 400 62130 430
rect 62246 400 62410 430
rect 62526 400 62690 430
rect 62806 400 62970 430
rect 63086 400 63250 430
rect 63366 400 63530 430
rect 63646 400 63810 430
rect 63926 400 64090 430
rect 64206 400 64370 430
rect 64486 400 64650 430
rect 64766 400 64930 430
rect 65046 400 65210 430
rect 65326 400 65490 430
rect 65606 400 65770 430
rect 65886 400 66050 430
rect 66166 400 66330 430
rect 66446 400 66610 430
rect 66726 400 66890 430
rect 67006 400 67170 430
rect 67286 400 67450 430
rect 67566 400 67730 430
rect 67846 400 68010 430
rect 68126 400 68290 430
rect 68406 400 68570 430
rect 68686 400 68850 430
rect 68966 400 69130 430
rect 69246 400 69410 430
rect 69526 400 69690 430
rect 69806 400 69970 430
rect 70086 400 70250 430
rect 70366 400 70530 430
rect 70646 400 70810 430
rect 70926 400 71090 430
rect 71206 400 71370 430
rect 71486 400 71650 430
rect 71766 400 71930 430
rect 72046 400 72210 430
rect 72326 400 72490 430
rect 72606 400 72770 430
rect 72886 400 73050 430
rect 73166 400 73330 430
rect 73446 400 73610 430
rect 73726 400 73890 430
rect 74006 400 74170 430
rect 74286 400 74450 430
rect 74566 400 74730 430
rect 74846 400 75010 430
rect 75126 400 75290 430
rect 75406 400 75570 430
rect 75686 400 75850 430
rect 75966 400 76130 430
rect 76246 400 76410 430
rect 76526 400 76690 430
rect 76806 400 76970 430
rect 77086 400 77250 430
rect 77366 400 77530 430
rect 77646 400 77810 430
rect 77926 400 78090 430
rect 78206 400 78370 430
rect 78486 400 78650 430
rect 78766 400 78930 430
rect 79046 400 79210 430
rect 79326 400 79490 430
rect 79606 400 79770 430
rect 79886 400 80050 430
rect 80166 400 80330 430
rect 80446 400 80610 430
rect 80726 400 80890 430
rect 81006 400 81170 430
rect 81286 400 81450 430
rect 81566 400 81730 430
rect 81846 400 82010 430
rect 82126 400 82290 430
rect 82406 400 82570 430
rect 82686 400 82850 430
rect 82966 400 83130 430
rect 83246 400 83410 430
rect 83526 400 83690 430
rect 83806 400 83970 430
rect 84086 400 84250 430
rect 84366 400 84530 430
rect 84646 400 84810 430
rect 84926 400 85090 430
rect 85206 400 85370 430
rect 85486 400 85650 430
rect 85766 400 85930 430
rect 86046 400 86210 430
rect 86326 400 86490 430
rect 86606 400 86770 430
rect 86886 400 87050 430
rect 87166 400 89306 430
<< obsm3 >>
rect 9 1246 89087 58422
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 4494 2921 9874 6599
rect 10094 2921 17554 6599
rect 17774 2921 25234 6599
rect 25454 2921 32914 6599
rect 33134 2921 40594 6599
rect 40814 2921 48274 6599
rect 48494 2921 55954 6599
rect 56174 2921 60074 6599
<< labels >>
rlabel metal2 s 672 59600 728 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24192 59600 24248 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 26544 59600 26600 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 28896 59600 28952 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 31248 59600 31304 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 33600 59600 33656 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 35952 59600 36008 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38304 59600 38360 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40656 59600 40712 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43008 59600 43064 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45360 59600 45416 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3024 59600 3080 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47712 59600 47768 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50064 59600 50120 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 52416 59600 52472 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 54768 59600 54824 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57120 59600 57176 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 59472 59600 59528 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 61824 59600 61880 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 64176 59600 64232 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 66528 59600 66584 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 68880 59600 68936 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5376 59600 5432 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 71232 59600 71288 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 73584 59600 73640 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 75936 59600 75992 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 78288 59600 78344 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 80640 59600 80696 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 82992 59600 83048 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 85344 59600 85400 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 87696 59600 87752 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7728 59600 7784 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10080 59600 10136 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12432 59600 12488 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14784 59600 14840 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17136 59600 17192 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19488 59600 19544 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 21840 59600 21896 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1456 59600 1512 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 24976 59600 25032 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27328 59600 27384 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29680 59600 29736 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32032 59600 32088 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34384 59600 34440 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36736 59600 36792 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39088 59600 39144 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41440 59600 41496 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 43792 59600 43848 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46144 59600 46200 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3808 59600 3864 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48496 59600 48552 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 50848 59600 50904 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 53200 59600 53256 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 55552 59600 55608 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 57904 59600 57960 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 60256 59600 60312 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 62608 59600 62664 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 64960 59600 65016 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 67312 59600 67368 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 69664 59600 69720 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6160 59600 6216 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 72016 59600 72072 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 74368 59600 74424 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 76720 59600 76776 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 79072 59600 79128 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 81424 59600 81480 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 83776 59600 83832 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 86128 59600 86184 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 88480 59600 88536 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8512 59600 8568 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10864 59600 10920 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13216 59600 13272 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15568 59600 15624 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17920 59600 17976 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20272 59600 20328 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 22624 59600 22680 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2240 59600 2296 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 25760 59600 25816 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28112 59600 28168 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 30464 59600 30520 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 32816 59600 32872 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35168 59600 35224 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 39872 59600 39928 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42224 59600 42280 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44576 59600 44632 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 46928 59600 46984 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4592 59600 4648 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 49280 59600 49336 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 51632 59600 51688 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 53984 59600 54040 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 56336 59600 56392 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 58688 59600 58744 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 61040 59600 61096 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 63392 59600 63448 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 65744 59600 65800 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 68096 59600 68152 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 70448 59600 70504 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6944 59600 7000 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 72800 59600 72856 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 75152 59600 75208 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 77504 59600 77560 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 79856 59600 79912 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 82208 59600 82264 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 84560 59600 84616 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 86912 59600 86968 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 89264 59600 89320 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9296 59600 9352 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11648 59600 11704 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14000 59600 14056 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16352 59600 16408 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18704 59600 18760 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 21056 59600 21112 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 86240 0 86296 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 86520 0 86576 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 86800 0 86856 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 32480 0 32536 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 41720 0 41776 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 42560 0 42616 400 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 43400 0 43456 400 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 45080 0 45136 400 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 46760 0 46816 400 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 48440 0 48496 400 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 33320 0 33376 400 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 49280 0 49336 400 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 50120 0 50176 400 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 51800 0 51856 400 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 53480 0 53536 400 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 55160 0 55216 400 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 56000 0 56056 400 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 56840 0 56896 400 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 57680 0 57736 400 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 58520 0 58576 400 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 60200 0 60256 400 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 61040 0 61096 400 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 61880 0 61936 400 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 62720 0 62776 400 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 63560 0 63616 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 64400 0 64456 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 65240 0 65296 400 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 35000 0 35056 400 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 66920 0 66976 400 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 67760 0 67816 400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 68600 0 68656 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 69440 0 69496 400 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 70280 0 70336 400 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 71120 0 71176 400 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 71960 0 72016 400 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 73640 0 73696 400 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 74480 0 74536 400 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 75320 0 75376 400 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 76160 0 76216 400 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 77000 0 77056 400 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 77840 0 77896 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 78680 0 78736 400 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 79520 0 79576 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 80360 0 80416 400 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 81200 0 81256 400 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 82040 0 82096 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 36680 0 36736 400 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 82880 0 82936 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 83720 0 83776 400 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 84560 0 84616 400 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 85400 0 85456 400 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 37520 0 37576 400 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 38360 0 38416 400 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 40040 0 40096 400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 32760 0 32816 400 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 41160 0 41216 400 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 42000 0 42056 400 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 42840 0 42896 400 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 43680 0 43736 400 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 44520 0 44576 400 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 46200 0 46256 400 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 47880 0 47936 400 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 48720 0 48776 400 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 33600 0 33656 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 49560 0 49616 400 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 51240 0 51296 400 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 52920 0 52976 400 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 54600 0 54656 400 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 55440 0 55496 400 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 56280 0 56336 400 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 34440 0 34496 400 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 57960 0 58016 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 58800 0 58856 400 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 59640 0 59696 400 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 60480 0 60536 400 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 61320 0 61376 400 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 62160 0 62216 400 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 63000 0 63056 400 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 63840 0 63896 400 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 64680 0 64736 400 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 65520 0 65576 400 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 35280 0 35336 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 66360 0 66416 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 67200 0 67256 400 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 68040 0 68096 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 68880 0 68936 400 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 69720 0 69776 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 70560 0 70616 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 71400 0 71456 400 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 72240 0 72296 400 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 73080 0 73136 400 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 73920 0 73976 400 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 36120 0 36176 400 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 74760 0 74816 400 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 75600 0 75656 400 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 76440 0 76496 400 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 77280 0 77336 400 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 78120 0 78176 400 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 78960 0 79016 400 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 79800 0 79856 400 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 80640 0 80696 400 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 81480 0 81536 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 82320 0 82376 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 36960 0 37016 400 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 83160 0 83216 400 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 84000 0 84056 400 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 84840 0 84896 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 85680 0 85736 400 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 37800 0 37856 400 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 39480 0 39536 400 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 40320 0 40376 400 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 33040 0 33096 400 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 42280 0 42336 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 43960 0 44016 400 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 44800 0 44856 400 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 45640 0 45696 400 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 46480 0 46536 400 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 47320 0 47376 400 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 49000 0 49056 400 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 33880 0 33936 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 50680 0 50736 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 51520 0 51576 400 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 52360 0 52416 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 54040 0 54096 400 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 55720 0 55776 400 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 56560 0 56616 400 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 57400 0 57456 400 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 58240 0 58296 400 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 59080 0 59136 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 60760 0 60816 400 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 62440 0 62496 400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 64120 0 64176 400 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 64960 0 65016 400 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 65800 0 65856 400 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 35560 0 35616 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 66640 0 66696 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 67480 0 67536 400 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 68320 0 68376 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 69160 0 69216 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 70000 0 70056 400 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 70840 0 70896 400 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 71680 0 71736 400 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 72520 0 72576 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 73360 0 73416 400 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 74200 0 74256 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 75040 0 75096 400 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 75880 0 75936 400 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 77560 0 77616 400 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 78400 0 78456 400 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 79240 0 79296 400 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 80080 0 80136 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 80920 0 80976 400 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 81760 0 81816 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 82600 0 82656 400 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 37240 0 37296 400 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 84280 0 84336 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 85120 0 85176 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 85960 0 86016 400 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 38080 0 38136 400 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 38920 0 38976 400 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 39760 0 39816 400 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 40600 0 40656 400 6 la_oenb[9]
port 309 nsew signal input
rlabel metal2 s 87080 0 87136 400 6 user_clock2
port 310 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 2800 0 2856 400 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 3080 0 3136 400 6 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 4480 0 4536 400 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 14840 0 14896 400 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 16520 0 16576 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 17360 0 17416 400 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 18200 0 18256 400 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 19880 0 19936 400 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 21560 0 21616 400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 22400 0 22456 400 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 23240 0 23296 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 24920 0 24976 400 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 26600 0 26656 400 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 28280 0 28336 400 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 29120 0 29176 400 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 29960 0 30016 400 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 31640 0 31696 400 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 9800 0 9856 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 11480 0 11536 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 12320 0 12376 400 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 13160 0 13216 400 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 3640 0 3696 400 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 4760 0 4816 400 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 14280 0 14336 400 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 15960 0 16016 400 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 17640 0 17696 400 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 19320 0 19376 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 21000 0 21056 400 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 5880 0 5936 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 22680 0 22736 400 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 24360 0 24416 400 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 26040 0 26096 400 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 27720 0 27776 400 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 29400 0 29456 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 7000 0 7056 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 31080 0 31136 400 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 8120 0 8176 400 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 9240 0 9296 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 10920 0 10976 400 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 12600 0 12656 400 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 14560 0 14616 400 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 15400 0 15456 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 17080 0 17136 400 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 17920 0 17976 400 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 18760 0 18816 400 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 20440 0 20496 400 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 21280 0 21336 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 22120 0 22176 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 6160 0 6216 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 22960 0 23016 400 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 23800 0 23856 400 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 24640 0 24696 400 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 25480 0 25536 400 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 26320 0 26376 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 27160 0 27216 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 28000 0 28056 400 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 28840 0 28896 400 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 30520 0 30576 400 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 7280 0 7336 400 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 31360 0 31416 400 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 32200 0 32256 400 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 9520 0 9576 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 10360 0 10416 400 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 11200 0 11256 400 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 12040 0 12096 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 12880 0 12936 400 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 13720 0 13776 400 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 5320 0 5376 400 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 6440 0 6496 400 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 7560 0 7616 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 8680 0 8736 400 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 3920 0 3976 400 6 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 4200 0 4256 400 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3704724
string GDS_FILE /home/passant/caravel_user_project-gf180mcu/openlane/user_proj_example/runs/22_12_11_11_17/results/signoff/user_proj_example.magic.gds
string GDS_START 78210
<< end >>

